<%
	proc writeTemplate {object} {
		
		$object onEachComponent {
			if {[$it isa osys::rfg::Group]} {
				writeTemplate $it
			} else {
				set register $it
				$it onEachField {
					puts "	.[$register name]_[$it name](),"				
				}
			}
		}

	}
	
	proc writeBlackbox {registerFile} {
		puts "writeBlackbox"
	}

	proc writeRegisternames {registerFile} {
		puts "writeRegisternames"
	}

	proc writeRegister {registerFile} {
		puts "writeRegister"
	}

	proc writeAddressControl {registerFile} {
		puts "writeAddressControl"
	}
%>
/* auto generated by RFG */
/*
<%puts -nonewline "[$registerFile name] [$registerFile name]"%>_I (
	.res_n(),
	.clk(),
	.address(),
	.read_data(),
	.invalid_address(),
	.access_complete(),
	.read_en(),
	.write_en(),
	.write_data(),
<% writeTemplate $registerFile %>);
*/
module <%puts [$registerFile name]%>(
	<% writeBlackbox $registerFile %>
);

<% writeRegisternames $registerFile %>

<% writeRegister $registerFile %>

<% writeAddressControl $registerFile %>

endmodule;